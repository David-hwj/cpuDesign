LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY zhiling IS
	PORT(
	EN		:IN STD_LOGIC;
	IRR		:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	MOVA	:OUT STD_LOGIC;
	MOVB	:OUT STD_LOGIC;
	MOVC	:OUT STD_LOGIC;
	ADD,SUB,AND0		:OUT STD_LOGIC;
	NOT0	:OUT STD_LOGIC;
	SHL		:OUT STD_LOGIC;
	SHR		:OUT STD_LOGIC;
	JZ,JC,IN0,OUT0,JMP,NOP:OUT STD_LOGIC;
	HALT	:OUT STD_LOGIC);
END zhiling;

ARCHITECTURE BEHAV OF zhiling IS
SIGNAL DATA		:STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN
	DATA <= IRR(7) & IRR(6) & IRR(5) & IRR(4);
	PROCESS(DATA,IRR)
	VARIABLE ZMOVA	:STD_LOGIC;
	VARIABLE ZMOVB	:STD_LOGIC;
	VARIABLE ZMOVC	:STD_LOGIC;
	VARIABLE ZADD,ZAND0,ZJZ,ZJC,ZIN0,ZOUT0,ZNOP,ZJMP,ZSUB	:STD_LOGIC;
	VARIABLE ZNOT0	:STD_LOGIC;
	VARIABLE ZSHL	:STD_LOGIC;
	VARIABLE ZSHR	:STD_LOGIC;
	VARIABLE ZHALT	:STD_LOGIC;
	BEGIN
	ZMOVA	:='0';
	ZMOVB	:='0';
	ZMOVC	:='0';
	ZADD	:='0';
	ZAND0	:='0';
	ZJZ		:='0';
	ZJC		:='0';
	ZIN0	:='0';
	ZOUT0   :='0';
	ZJMP	:='0';
	ZNOP	:='0';
	ZSUB	:='0';
	ZNOT0	:='0';
	ZSHL	:='0';
	ZSHR	:='0';
	ZHALT	:='0';
			IF(DATA = "0011") THEN
				IF(IRR(3 DOWNTO 2) = "11") THEN
					ZMOVB:='1';	
				ELSIF(IRR(1 DOWNTO 0) = "11") THEN
					ZMOVC:='1';
				ELSE
					ZMOVA:='1';
				END IF;
			ELSIF(DATA = "1001") THEN
				ZADD:='1';
			ELSIF(DATA = "0110") THEN
				ZSUB:='1';
			ELSIF(DATA = "1110") THEN
				ZAND0:='1';
			ELSIF(DATA = "0101") THEN
				ZNOT0:='1';
			ELSIF(DATA = "0010") THEN
				ZIN0:='1';
			ELSIF(DATA = "0100") THEN
				ZOUT0:='1';
			ELSIF(DATA = "1010") THEN
				IF(IRR(1 DOWNTO 0) = "00") THEN
					ZSHR:='1';
				ELSIF(IRR(1 DOWNTO 0) = "11") THEN
					ZSHL:='1';
				END IF;
			ELSIF IRR="10000000" THEN
				ZHALT:='1';
			ELSIF(DATA = "0001") THEN
				IF(IRR(1 DOWNTO 0) = "00") THEN
					ZJMP:='1';
				ELSIF(IRR(1 DOWNTO 0) = "01") THEN
					ZJZ:='1';				
				ELSIF(IRR(1 DOWNTO 0) = "10") THEN
					ZJC:='1';
				END IF;
			END IF;
			IF(EN='0')THEN
	ZMOVA	:='0';
	ZMOVB	:='0';
	ZMOVC	:='0';
	ZADD	:='0';
	ZAND0	:='0';
	ZJZ		:='0';
	ZJC		:='0';
	ZIN0	:='0';
	ZOUT0   :='0';
	ZJMP	:='0';
	ZNOP	:='0';
	ZSUB	:='0';
	ZNOT0	:='0';
	ZSHL	:='0';
	ZSHR	:='0';
	ZHALT	:='0';
			END IF;
			MOVA<=ZMOVA;
			MOVB<=ZMOVB;
			MOVC<=ZMOVC;
			ADD<=ZADD;
			SUB<=ZSUB;
			AND0<=ZAND0;
			JZ<=ZJZ;
			JC<=ZJC;
			IN0<=ZIN0;
			OUT0<=ZOUT0;
			JMP<=ZJMP;
			NOP<=ZNOP;
			NOT0<=ZNOT0;
			SHL<=ZSHL;
			SHR<=ZSHR;
			HALT<=ZHALT;
	END PROCESS;
END BEHAV;
