lpm_decode0_inst : lpm_decode0 PORT MAP (
		data	 => data_sig,
		eq3	 => eq3_sig
	);
